interface dut_if();
  logic clk;
  logic rst_n;
endinterface