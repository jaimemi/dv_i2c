`include "base_test.sv"

`include "test_dummy.sv"
//other tests
`include "test_write.sv"
`include "test_read.sv"
`include "test_rw_rand.sv"
`include "test_clk.sv"
`include "test_abort.sv"
`include "test_device_addr.sv"
`include "test_all.sv"