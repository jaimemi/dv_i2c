`include "base_test.sv"

`include "test_dummy.sv"
//other tests
`include "test_write.sv"